`include "apb_interface.sv"
`include "top.sv"
