`ifndef APB_TEST_PKG
`define APB_TEST_PKG

package apb_test_pkg;
  import uvm_pkg::*
  `include "uvm_macros.svh";
  
  import apb_agent_pkg::*;
  import apb_sequence_pkg::*;
  import apb_env_pkg::*;

  `include "apb_test_cfg.sv"
  `include "apb_base_test.sv"
  `include "apb_valid_rw_test.sv"
  `include "apb_err_rw_test.sv"
  `include "apb_mem_integrity_test.sv"
  `include "apb_rand_test.sv"
endpackage
`endif
