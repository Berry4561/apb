`ifndef APB_ENV_PKG
`define APB_ENV_PKG

package apb_env_pkg;
  import uvm_pkg::*
  `include "uvm_macros.svh";

  import apb_agent_pkg::*;

  `include "apb_dut_checker.sv"
  `include "apb_env.sv"
endpackage
`endif
