`include "apb_interface.sv"
`include "apb_agent_pkg.sv"
`include "apb_sequence_pkg.sv"
`include "apb_env_pkg.sv"
`include "apb_test_pkg.sv"

`include "top.sv"
