//THis file is the top module of the Testbench

module top;

endmodule
