`ifndef APB_SEQUENCE_PKG
`define APB_SEQUENCE_PKG

package apb_sequence_pkg;
  
  import uvm_pkg::*;
  `include "uvm_macros.svh";

  import apb_agent_pkg::*;
  `include "apb_sequence.sv"

endpackage
`endif
