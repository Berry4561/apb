`ifndef APB_AGENT_PKG
`define APB_AGENT_PKG

package apb_agent_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "apb_transaction.sv"
  `include "apb_sequence.sv"
  `include "apb_sequnecer.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  `include "apb_agent.sv"
endpackage
`endif
