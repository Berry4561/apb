//THis file is the top module of the Testbench

module top;

  //apb_interface apb_if();
  
  //apb_dut dut1();

  //CLock GEN Block;
  
endmodule
