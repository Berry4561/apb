`include "apb_top.sv";
